module downcounter_testbench();
reg clk, reset;
wire [3:0] counter;
down_counter dut(clk, reset, counter);
initial begin 
clk=0;
forever #5 clk=~clk;
end
initial begin
		$dumpfile("dump.vcd");
			$dumpvars(0,downcounter_testbench);
reset=1;
#20;
reset=0;
end
endmodule 
