 //Module magnitude comparator 
module magnitude_comparator(A_gt_B, A_lt_B, A_eq_B, A, B); 
//Comparison output 
output A_gt_B, A_lt_B, A_eq_B; 
//4-bits numbers input 
input [3:0] A, B; 
assign A_gt_B = (A > B); //A greater than B 
assign A_lt_B = (A < B); //A less than B 
assign A_eq_B = (A == B); //A equal to B 
endmodule
